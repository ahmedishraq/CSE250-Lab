* H:\Circuit Design\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Mon Nov 01 20:12:31 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
